// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
module mac_tile (clk, out_s, in_w, out_e, in_n, inst_w, inst_e, reset);
parameter bw = 4;
parameter psum_bw = 16;

output [psum_bw-1:0] out_s;
input  [bw-1:0] in_w; 
output [bw-1:0] out_e; 
input  [2:0] inst_w; 
//inst[2] == 1: output_stationary, inst[1]:pass_psum, inst[0]: accumulate
//inst[2] == 0: weight stationary, inst[1]:execute, inst[0]: kernel loading
output [2:0] inst_e;
input  [psum_bw-1:0] in_n;  //either weight from output_stationary or psum from weight stationary
input  clk;
input  reset;
wire weight_stationary;
assign weight_stationary = ~inst[2];
reg [bw-1:0] a_q
reg [psum_bw-1:0] b_q;
reg [psum_bw-1:0] c_q;
reg [1:0] inst_q;
reg load_ready_q;

wire signed [psum_bw-1:0] mac_out; 
mac #(.bw(bw), .psum_bw(psum_bw)) mac_instance (
    .a(a_q), 
    .b(b_q),
    .c(c_q),
    .out(mac_out)
); 
always @(posedge clk) begin
    if (reset) begin
        inst_q <= 2'b00;
        load_ready_q <= 1;
        a_q <= 0;
        b_q <= 0;
        c_q <= 0;

    end else if (weight_stationary) begin    //weight stationary
        inst_q[1] <= inst_w[1]; // Accept your inst_w[1] (execution) always into inst_q[1] latch.
        if (inst_w[1] == 1 || inst_w[0] == 1) begin
            a_q <= in_w;
        end

        if (inst_w[0] == 1 && load_ready_q == 1) begin
            b_q <= in_w; // b_q holds the weights
            load_ready_q <= 0;
        end

        c_q <= in_n;
        
        if (load_ready_q == 0) begin
            inst_q[0] <= inst_w[0];
        end
    end else begin  //output stationary
        inst_q = inst_w; // Question: should the instructions be passed down no matter what? Yes? Yes.
        if(inst_w[0]) begin//inst[2] == 1: output_stationary, inst[1]:pass_psum, inst[0]: accumulate
        a_q = in_w;
        b_q = in_n;
        end

    end 
end

//In output stationary case, we need to get mac_out into c_q before next posedge
//(a_q and b_q will be changed at next rising edge and thus changing mac_out).
always @ (negedge clk) begin
    if(inst_w[0] && inst_w[2]) begin
        c_q = mac_out
    end
end

assign out_e = a_q;
assign inst_e = inst_q;
assign out_s = inst[2] ? (inst [1] ? c_q : b_q) :mac_out; // if output stationary, pass down weight. Else, pass down psum
endmodule
