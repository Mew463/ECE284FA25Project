// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module mac_row (clk, out_s, in_w, in_n, valid, inst_w, reset, weight_stationary, pass_psum, recall_psum);

  parameter bw = 4;
  parameter psum_bw = 16;
  parameter col = 8;

  input  clk, reset;
  output [psum_bw*col-1:0] out_s;
  output [col-1:0] valid;
  // inst[1]:execute, inst[0]: kernel loading
  input  [bw-1:0] in_w; 
  input  [1:0] inst_w; 
  input  [psum_bw*col-1:0] in_n;
  input pass_psum, weight_stationary, recall_psum;

  wire  [(col+1)*bw-1:0] temp; // Temp is passing either weights or the input
  wire  [(col+1)*2:0] inst_temp; // Passing instruction

  assign temp[bw-1:0]   = in_w;
  assign inst_temp[1:0] = inst_w;

  genvar i;
  for (i=1; i < col+1 ; i=i+1) begin : col_num
      mac_tile #(.bw(bw), .psum_bw(psum_bw)) mac_tile_instance (
        .clk(clk),
        .reset(reset),
        .in_w( temp[bw*(i-1)+: bw]),
        .out_e(temp[bw*i +: bw]),
        .inst_w(inst_temp[2*(i-1) +: 2]),
        .inst_e(inst_temp[2*i +: 2]),
        .in_n(in_n[psum_bw*(i-1) +: psum_bw]),
        .out_s(out_s[psum_bw*(i-1) +: psum_bw]),
        .weight_stationary(weight_stationary),
        .pass_psum(pass_psum),
        .recall_psum(recall_psum));

   assign valid[i-1] = inst_temp[2*i+1]; // " valid for the column is inst_e[1] for the column"
  end

endmodule
