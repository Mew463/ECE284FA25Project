module core;

parameter bw = 4;
parameter psum_bw = 16;
